package CodicInterface;

import ClientServer :: *;
import FloatingPoint :: *;


typedef Server  #(Float) CordicIFC;


endpackage
