// e^x using CORDIC Alogrithm 