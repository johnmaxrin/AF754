package CordicInterface;

import ClientServer :: *;
import FloatingPoint :: *;

interface CordicIFC;
    interface Server  #(Bit#(16), Bit#(16)) cordicServerIFC;
    //method Action dometh(Bit#(16));
endinterface

endpackage
